  
  `define READ_ROM  8'h33
  `define MATCH_ROM  8'h55

  `define READ_SCRPD  8'h3e
  `define WRITE_SCRPD 8'hbe
  
  `define UID_DATA 56'h98765432109876
  
  
  
 
