module ows_wr_interface (
	input clk,
	input snd_prsnc,
	
	output data_out,
	output data_out_oe
);

endmodule
